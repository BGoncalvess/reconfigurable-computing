library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


entity noisy_signal is
    Port ( 
        addr : in unsigned(9 downto 0);
        data_out : out signed(15 downto 0)
    );
end noisy_signal;

architecture Behaviroal of noisy_signal is 

    
type signal_value is array (0 to 999) of signed(15 downto 0);

-- Declare the constant using the defined type
constant signal_array : signal_value := (
    signed(1111111110100010),
    signed(1111101010110000),
    signed(0000101100001111),
    signed(0001100101000010),
    signed(0001011000100101),
    signed(0010101010100010),
    signed(0010001000110011),
    signed(0010111110101100),
    signed(0011010101101000),
    signed(0100011110011011),
    signed(0011110111010100),
    signed(0011101100100000),
    signed(0011100110101010),
    signed(0100111001111001),
    signed(0100010101100011),
    signed(0101011111100000),
    signed(0100110100011011),
    signed(0100011001111100),
    signed(0011111111101000),
    signed(0100000001110011),
    signed(0011101101010011),
    signed(0011110100000110),
    signed(0011111000010101),
    signed(0100110000100101),
    signed(0011001111110110),
    signed(0100001101100110),
    signed(0011101111001110),
    signed(0101001010110000),
    signed(0100100000101110),
    signed(0100001001011111),
    signed(0011111010011111),
    signed(0101000110000100),
    signed(0100001111110101),
    signed(0110011110001000),
    signed(0101000010011110),
    signed(0100010000100001),
    signed(0101011011110101),
    signed(0101110101101001),
    signed(0101111000000110),
    signed(0101000000110001),
    signed(0011110011001010),
    signed(0100000100011110),
    signed(0100101011110100),
    signed(0100001100101010),
    signed(0100001100000100),
    signed(0100000101001001),
    signed(0011110110111010),
    signed(0011010110100101),
    signed(0011101011000101),
    signed(0011011011101010),
    signed(0001110011110100),
    signed(0010000000010000),
    signed(0001101010001111),
    signed(0010110101111100),
    signed(0000111101101111),
    signed(0000110111111100),
    signed(0000100010101100),
    signed(1111110001011011),
    signed(1111010001000011),
    signed(1111111001100101),
    signed(0000001100001010),
    signed(0000111011110011),
    signed(0000010001010110),
    signed(0000001100100011),
    signed(0000101000011110),
    signed(0000011011010101),
    signed(0000101110010100),
    signed(1111111000100001),
    signed(0001010111111000),
    signed(0010000001011011),
    signed(0001110110100001),
    signed(0010011111011111),
    signed(0001010001000011),
    signed(0010001000110101),
    signed(0001010001100000),
    signed(0001111000111110),
    signed(0001101000100001),
    signed(0001100101101111),
    signed(0010011111111111),
    signed(0001110011000110),
    signed(0010100001111100),
    signed(0011111011111100),
    signed(0001010110000111),
    signed(0010100010010011),
    signed(0010000111001010),
    signed(0001110001011000),
    signed(0010011110100111),
    signed(0001001000100011),
    signed(0001010101111100),
    signed(0000111111000101),
    signed(0001110100110111),
    signed(0000010111011100),
    signed(0000001110011111),
    signed(0001011101100111),
    signed(0001001000011000),
    signed(0001110100010000),
    signed(0001011111101100),
    signed(0001100111111000),
    signed(0001111110110000),
    signed(0001001011011001),
    signed(0010011000101111),
    signed(0010110000011100),
    signed(0010101011110011),
    signed(0011100100011100),
    signed(0011000111001110),
    signed(0010111111100011),
    signed(0011101100010001),
    signed(0011001100001000),
    signed(0010110110101011),
    signed(0010001000001110),
    signed(0010101010000010),
    signed(0001110101111100),
    signed(0001000100011010),
    signed(0001100110010111),
    signed(0000101100110001),
    signed(0000101010100111),
    signed(1111010111011011),
    signed(0000001010111100),
    signed(1110011111111000),
    signed(1110100001011111),
    signed(1110000011011111),
    signed(1110101101110110),
    signed(1110001001110011),
    signed(1101100101100010),
    signed(1100010101001000),
    signed(1011001000011011),
    signed(1011001101000100),
    signed(1100010010110101),
    signed(1011111000000110),
    signed(1100111101000110),
    signed(1001110011000000),
    signed(1011011010010011),
    signed(1010101100110010),
    signed(1100101011110010),
    signed(1011011111111101),
    signed(1100001101000001),
    signed(1011010000001101),
    signed(1011011111110000),
    signed(1011111001111001),
    signed(1100000110101001),
    signed(1011101101010010),
    signed(1010011011101100),
    signed(1011011101000101),
    signed(1010011110111001),
    signed(1010111001001010),
    signed(1010110010000010),
    signed(1010000100101000),
    signed(1011011100101111),
    signed(1010100000000110),
    signed(1010010010011011),
    signed(1001010010110001),
    signed(1001110000101001),
    signed(1000011010111111),
    signed(1001101011111101),
    signed(1001000001110100),
    signed(1001010001000110),
    signed(1010000010001001),
    signed(1000000101000010),
    signed(1010010100101000),
    signed(1010100001100110),
    signed(1001101101011111),
    signed(1010001100101010),
    signed(1100000010001011),
    signed(1011100111010010),
    signed(1010111101111010),
    signed(1011000101110111),
    signed(1101001000111100),
    signed(1100010011101011),
    signed(1101100011110101),
    signed(1110010000001011),
    signed(1110100000110001),
    signed(1110100001110111),
    signed(1111110111001001),
    signed(1111110001101010),
    signed(1110101000000101),
    signed(1111110011010100),
    signed(1111110010111111),
    signed(0000111010110110),
    signed(0001100000000011),
    signed(0000010101000100),
    signed(0000100100001111),
    signed(0000110100001010),
    signed(1111111110100010),
    signed(1111001111101111),
    signed(1111111010000010),
    signed(0000101010110110),
    signed(0000101000100110),
    signed(0000101100010110),
    signed(0000001011001010),
    signed(0000011100101101),
    signed(1111010001001000),
    signed(1111100110010111),
    signed(0000101001011000),
    signed(1111111011100000),
    signed(0000110011010011),
    signed(0000011110100001),
    signed(0000100101100111),
    signed(0000111111010010),
    signed(0001101111010000),
    signed(0000010001101100),
    signed(0001101100110110),
    signed(0010000000111001),
    signed(0010000100110111),
    signed(0010100110110101),
    signed(0001111110011100),
    signed(0010001010110010),
    signed(0010010100000000),
    signed(0010000000000111),
    signed(0001111101011000),
    signed(0001101110010101),
    signed(0010000110010011),
    signed(0001100001111011),
    signed(0001001110110000),
    signed(0001110001010011),
    signed(0001001001111000),
    signed(0010100011011001),
    signed(1111111000001100),
    signed(0000001111100001),
    signed(0001001001011110),
    signed(1111001110110101),
    signed(1111011100011010),
    signed(1111001110000001),
    signed(1111010101100000),
    signed(1110101101000010),
    signed(1111000010101101),
    signed(1110101110100001),
    signed(1111010110100111),
    signed(1110110011011000),
    signed(1110101110101000),
    signed(0000000110100001),
    signed(1111111111011100),
    signed(0000111111000111),
    signed(0001001100001110),
    signed(0000111000010011),
    signed(0010001011111011),
    signed(0001111011101101),
    signed(0001101001111110),
    signed(0010010111000011),
    signed(0010010010011101),
    signed(0010010001100000),
    signed(0011111000001101),
    signed(0011101010000101),
    signed(0100010100110010),
    signed(0011000010100010),
    signed(0011101011110000),
    signed(0011110000011111),
    signed(0011010111001011),
    signed(0011101000101101),
    signed(0011100101100110),
    signed(0011011000100110),
    signed(0011100110010000),
    signed(0011001011111110),
    signed(0100001001011000),
    signed(0011001001100011),
    signed(0011000111001101),
    signed(0100100110111100),
    signed(0011001001010111),
    signed(0011010010001111),
    signed(0011011111110110),
    signed(0011010001110101),
    signed(0100100001110111),
    signed(0100100011101100),
    signed(0100000000110100),
    signed(0101001010001001),
    signed(0101001101111110),
    signed(0101001011100111),
    signed(0100011110101101),
    signed(0100101000101100),
    signed(0110011110110110),
    signed(0110010011001110),
    signed(0101110111110000),
    signed(0101111001001001),
    signed(0101110111111000),
    signed(0111100100010010),
    signed(0110010100111101),
    signed(0110000111101010),
    signed(0101101100011000),
    signed(0101111100011110),
    signed(0110110010101010),
    signed(0101001010101000),
    signed(0100110000111000),
    signed(0011111101101011),
    signed(0100010001111100),
    signed(0010110010001001),
    signed(0010010110101111),
    signed(0010000100010111),
    signed(0010010000010111),
    signed(0001101110100011),
    signed(0000111111000110),
    signed(0000011001001011),
    signed(1111110101010010),
    signed(1111111101010111),
    signed(0000000111101111),
    signed(1111001010100001),
    signed(0000000001110100),
    signed(1110101100100000),
    signed(1110101101100110),
    signed(1110100111101000),
    signed(1110011010110011),
    signed(1110011001000101),
    signed(1110100111101010),
    signed(1110000011001011),
    signed(1110010111001100),
    signed(1110111000100101),
    signed(1101111000010110),
    signed(1101111110101000),
    signed(1110010011111010),
    signed(1101101101010001),
    signed(1110000001001100),
    signed(1101000100111010),
    signed(1100110110110111),
    signed(1100101101000100),
    signed(1101011001100111),
    signed(1100111101100000),
    signed(1100111010011110),
    signed(1100010110101011),
    signed(1101000100001010),
    signed(1100011101001100),
    signed(1011110001000110),
    signed(1011100111001110),
    signed(1011010111101111),
    signed(1010011111011110),
    signed(1010111010110001),
    signed(1010110101001000),
    signed(1011110011111110),
    signed(1011100101101111),
    signed(1010100101011000),
    signed(1010100100001001),
    signed(1010110010001101),
    signed(1011100101001110),
    signed(1100100000110000),
    signed(1100101000000010),
    signed(1100111010011000),
    signed(1101010110011111),
    signed(1100001111011101),
    signed(1101000011000111),
    signed(1101101111111000),
    signed(1101111110000111),
    signed(1110010101001001),
    signed(1111000111000001),
    signed(1110101100001110),
    signed(1110100010111001),
    signed(1111101100000011),
    signed(1110111011101100),
    signed(1111001111110100),
    signed(1110110101000011),
    signed(1101110111010110),
    signed(1110100001111011),
    signed(1111000000000010),
    signed(1110011010010110),
    signed(1101110111111100),
    signed(1100110101000001),
    signed(1111010100111011),
    signed(1110000110111101),
    signed(1110010000001001),
    signed(1110010011011111),
    signed(1100100110000110),
    signed(1101010111011001),
    signed(1110000100011100),
    signed(1101001001101111),
    signed(1101110101010100),
    signed(1110101110001010),
    signed(1101111010100100),
    signed(1101101010000100),
    signed(1101101010100000),
    signed(1110001101010010),
    signed(1110101101111101),
    signed(1110111100111010),
    signed(1110000000001000),
    signed(0000000011100011),
    signed(1110101000111101),
    signed(1111010001010000),
    signed(1110100110111101),
    signed(1110101111001111),
    signed(1111000000000010),
    signed(1110111011110001),
    signed(1110000111101000),
    signed(1101001100101010),
    signed(1110110101001000),
    signed(1101101100100100),
    signed(1110000000011010),
    signed(1100111111110000),
    signed(1100011010110010),
    signed(1101011101111011),
    signed(1100100111010010),
    signed(1010011101001001),
    signed(1100000110100010),
    signed(1100001010110000),
    signed(1100000010011011),
    signed(1011110101101010),
    signed(1011100011001111),
    signed(1010111010100111),
    signed(1011111000110100),
    signed(1011001000101010),
    signed(1011110011010110),
    signed(1011100001011000),
    signed(1101000111000100),
    signed(1101001101111011),
    signed(1100010010101000),
    signed(1101100100101110),
    signed(1101001101111101),
    signed(1110110100011001),
    signed(1110111110100101),
    signed(1110111001001010),
    signed(1111101110011111),
    signed(1111100101011011),
    signed(1111000010100001),
    signed(0000001101011010),
    signed(0000001100111100),
    signed(0001010011001001),
    signed(0001011111001101),
    signed(0001010001011010),
    signed(0001110111110010),
    signed(0010011101101110),
    signed(0001000001001010),
    signed(0001011011111010),
    signed(0001011011111001),
    signed(0010000000011100),
    signed(0010011010010000),
    signed(0010110000101110),
    signed(0010011101001001),
    signed(0000000100111110),
    signed(0011010010111101),
    signed(0001001010110011),
    signed(0001101010110010),
    signed(0010110011011101),
    signed(0010101110100101),
    signed(0011101010001000),
    signed(0011011000101001),
    signed(0100001100011101),
    signed(0100101110011101),
    signed(0011000101100000),
    signed(0100101001101010),
    signed(0100111010001111),
    signed(0110010010000100),
    signed(0110001010101001),
    signed(0110000101111010),
    signed(0110101100001010),
    signed(0110101111010010),
    signed(0111111111111111),
    signed(0110111110000110),
    signed(0110101111011010),
    signed(0110110101100101),
    signed(0110110010000101),
    signed(0111011110100000),
    signed(0110110101010111),
    signed(0111110100000010),
    signed(0101110100111110),
    signed(0101101011000111),
    signed(0110100110110011),
    signed(0101111110100100),
    signed(0101010001001111),
    signed(0010111011011111),
    signed(0011000101001000),
    signed(0011001010110001),
    signed(0010100001011001),
    signed(0010001100101101),
    signed(0010000100110000),
    signed(0011101001101001),
    signed(0001111111101011),
    signed(0011000001011001),
    signed(0010001100111010),
    signed(0001011101001100),
    signed(0001011100111101),
    signed(0001111101111101),
    signed(0001101011110100),
    signed(0010011001100101),
    signed(0001001001010100),
    signed(0001111101100010),
    signed(0001100011101101),
    signed(0001001101100101),
    signed(0001001001001100),
    signed(0010001000000110),
    signed(0010000000101110),
    signed(0000110101100110),
    signed(0010011000111110),
    signed(0010011000000010),
    signed(0001010001000101),
    signed(1111010110010100),
    signed(0000000000000010),
    signed(0001100011010111),
    signed(0000011011011001),
    signed(0001010111011010),
    signed(1111110100010000),
    signed(1111101101001101),
    signed(1110100100110110),
    signed(1110010111001000),
    signed(1101001010010101),
    signed(1111001000101100),
    signed(1110001011000110),
    signed(1110011100111110),
    signed(1110101001101011),
    signed(1110111000111101),
    signed(1110011001101110),
    signed(1101111010111011),
    signed(1111001100001011),
    signed(1110010101101010),
    signed(1110011110001111),
    signed(1110101100010111),
    signed(1111110001101010),
    signed(1111111011000010),
    signed(0000010111111111),
    signed(0000011110111010),
    signed(0000101001100110),
    signed(0000110001001000),
    signed(0001101110101111),
    signed(0001100111110111),
    signed(0010011110000100),
    signed(0010101000100001),
    signed(0001110111111101),
    signed(0010001010111101),
    signed(0001100111110110),
    signed(0010101011011001),
    signed(0001101000010011),
    signed(0001001001010110),
    signed(0001100111111000),
    signed(0001011010110100),
    signed(0000011000010110),
    signed(0001001101011011),
    signed(0000000101001000),
    signed(1110101010000100),
    signed(1111000001010101),
    signed(1110010010101110),
    signed(1110101100011000),
    signed(1111001011001101),
    signed(1110001110000000),
    signed(1110111010110001),
    signed(1101111111011110),
    signed(1110100111111010),
    signed(1110000110111100),
    signed(1101101101110111),
    signed(1101110001011111),
    signed(1101110101011101),
    signed(1110111010111010),
    signed(1101110111011101),
    signed(1110110100011010),
    signed(1110000011011101),
    signed(1110000010011100),
    signed(1101011100000111),
    signed(1110011111010110),
    signed(1110100001100101),
    signed(1101000100010111),
    signed(1101000111110101),
    signed(1101101000100011),
    signed(1101010001001111),
    signed(1100101011111001),
    signed(1100110010110011),
    signed(1100001101000101),
    signed(1011100010011110),
    signed(1010000101001001),
    signed(1010101000001110),
    signed(1010101001010011),
    signed(1001001110001011),
    signed(1000111010010100),
    signed(1000111101001110),
    signed(1001000110101110),
    signed(1001101001000101),
    signed(1000110101101010),
    signed(1000100000001111),
    signed(1001101101001001),
    signed(1000111110001001),
    signed(1001101001001111),
    signed(1001110101110111),
    signed(1001011101100001),
    signed(1001001110111000),
    signed(1010010000100111),
    signed(1001111010010010),
    signed(1010001110011111),
    signed(1011000010011010),
    signed(1010110101101010),
    signed(1011100100011000),
    signed(1011111111100110),
    signed(1011110001001010),
    signed(1100101111011001),
    signed(1101001000000101),
    signed(1101100111101010),
    signed(1101111001001011),
    signed(1100111111001011),
    signed(1110010010111011),
    signed(1110010000000011),
    signed(1101110000010010),
    signed(1110100100001000),
    signed(1101101101011100),
    signed(1100001100110110),
    signed(1110011101010101),
    signed(1101111011001001),
    signed(1110000001000101),
    signed(1110111000001110),
    signed(1100111111010111),
    signed(1111001111101001),
    signed(1110011011110101),
    signed(0000001010101111),
    signed(1111000001011100),
    signed(1111011110101111),
    signed(0000010101000010),
    signed(0001000110100110),
    signed(0001010111111011),
    signed(0001100111110010),
    signed(0001011110101001),
    signed(0001110110111111),
    signed(0010001100001111),
    signed(0010111101110000),
    signed(0011000101111000),
    signed(0010110010110011),
    signed(0100000110001010),
    signed(0100101011001011),
    signed(0100001111001001),
    signed(0011111101111000),
    signed(0100010001000111),
    signed(0100101101101101),
    signed(0100101001011011),
    signed(0011101101110010),
    signed(0100111110101100),
    signed(0100100010111100),
    signed(0100010101111010),
    signed(0011101101110110),
    signed(0011111000101011),
    signed(0101001011100000),
    signed(0011001000010010),
    signed(0010010011010011),
    signed(0001000101100101),
    signed(0010010011111001),
    signed(0000101100011110),
    signed(0010101100010010),
    signed(0001111000101110),
    signed(0011010100111101),
    signed(0001100101010011),
    signed(0001010100111110),
    signed(0001111011010110),
    signed(0001111010011110),
    signed(0010000010110011),
    signed(0010000111000010),
    signed(0010011111000101),
    signed(0010000101001011),
    signed(0001101101011011),
    signed(0001101111010011),
    signed(0011000011010010),
    signed(0010011101101011),
    signed(0010110101010011),
    signed(0011001111111001),
    signed(0010001011011001),
    signed(0011001011000100),
    signed(0010101110101111),
    signed(0010010111001010),
    signed(0010101101100001),
    signed(0001000111010010),
    signed(0010101100000100),
    signed(0010100110000110),
    signed(0001001010001000),
    signed(0010100010000100),
    signed(0000100001101110),
    signed(0000100001011110),
    signed(1111111010010100),
    signed(0001110101110001),
    signed(1111111001101000),
    signed(0000100100001000),
    signed(0001000011011000),
    signed(0000100111011011),
    signed(0000001001101110),
    signed(0001001001101101),
    signed(0001100000010110),
    signed(0001110101110101),
    signed(0010000111101000),
    signed(0010011000010100),
    signed(0001101000111110),
    signed(0010111100001101),
    signed(0011100000011011),
    signed(0011001101110011),
    signed(0010111010011010),
    signed(0011110111011101),
    signed(0011011000101111),
    signed(0100110110011011),
    signed(0100010111100110),
    signed(0110010011001010),
    signed(0100100010101111),
    signed(0100101101011011),
    signed(0101010110011110),
    signed(0101111100101100),
    signed(0101010110110010),
    signed(0101110100010000),
    signed(0101111100101111),
    signed(0101000001111010),
    signed(0100101111101110),
    signed(0100000000101011),
    signed(0011110011001110),
    signed(0011100100111110),
    signed(0011011101101111),
    signed(0011100000011010),
    signed(0011111011110000),
    signed(0011100001110101),
    signed(0010001110111110),
    signed(0001010011000011),
    signed(0010010001010011),
    signed(0000101010000111),
    signed(0001011000101010),
    signed(0010100100101110),
    signed(0000101110010110),
    signed(0001010110001111),
    signed(0001000100111111),
    signed(0000111000111111),
    signed(0001010010010110),
    signed(0001011011000111),
    signed(0001001001011101),
    signed(0010000111110111),
    signed(0010000011000110),
    signed(0010110001001000),
    signed(0000100000010011),
    signed(1111010110000001),
    signed(0001001010101111),
    signed(1111101010100100),
    signed(1110111001111101),
    signed(1111010100111110),
    signed(1111100010000010),
    signed(1110111011101000),
    signed(1110111010111101),
    signed(1101001001001101),
    signed(1101010010100111),
    signed(1011111111011100),
    signed(1011001011100001),
    signed(1011011101011111),
    signed(1011000011100000),
    signed(1010100101011111),
    signed(1011110001111000),
    signed(1010011111011010),
    signed(1001111101101010),
    signed(1001101010010110),
    signed(1001101110100001),
    signed(1001110000010100),
    signed(1010010000000001),
    signed(1001111001110111),
    signed(1001010011101100),
    signed(1001110111100000),
    signed(1010010000010001),
    signed(1001010000100101),
    signed(1010000000010010),
    signed(1010110000100011),
    signed(1011001111111001),
    signed(1011111100110000),
    signed(1100000011010011),
    signed(1101001001111110),
    signed(1010010000001100),
    signed(1101000000001110),
    signed(1100010000101010),
    signed(1100010101111001),
    signed(1011110110111101),
    signed(1100100001100001),
    signed(1100111111101010),
    signed(1101010010111101),
    signed(1100111101110011),
    signed(1011110000001010),
    signed(1100001110100001),
    signed(1101000110011011),
    signed(1100001110010111),
    signed(1100000111110101),
    signed(1101010101011001),
    signed(1101011010010001),
    signed(1011011100001111),
    signed(1100011100100111),
    signed(1101010011011011),
    signed(1100001101111111),
    signed(1101010100111000),
    signed(1101100111000100),
    signed(1101101110100111),
    signed(1101111001000111),
    signed(1111011010111000),
    signed(1110100011101000),
    signed(1111010110100001),
    signed(0000001010000001),
    signed(1111000001110111),
    signed(1111100011010100),
    signed(1111111001111100),
    signed(0001010101110111),
    signed(0000111101000100),
    signed(0000101000001011),
    signed(0000001101101000),
    signed(0000010000101000),
    signed(0001101101100101),
    signed(0000000110001111),
    signed(0000001110101001),
    signed(0000111010111100),
    signed(1111110110011010),
    signed(0000011110001100),
    signed(1111101001001101),
    signed(1111110111111110),
    signed(1111010011000011),
    signed(1111011110100001),
    signed(1111100100100001),
    signed(1110111101101101),
    signed(1110010000100010),
    signed(1110111010011011),
    signed(1110001111011100),
    signed(1101001111000000),
    signed(1100100000100101),
    signed(1101110010001101),
    signed(1101010110101101),
    signed(1101101100111011),
    signed(1101010111001000),
    signed(1111010100010010),
    signed(1110001001110101),
    signed(1110101111110100),
    signed(1110001110010110),
    signed(1110110000111000),
    signed(1111111010010001),
    signed(1110101001011110),
    signed(1110101111000010),
    signed(1111011100011011),
    signed(0000011001111111),
    signed(0000100101001011),
    signed(1110010110001110),
    signed(1111100101101001),
    signed(1111110000000001),
    signed(0000100000101001),
    signed(0000100111010111),
    signed(1110100010111101),
    signed(1111011111111001),
    signed(1111110001011111),
    signed(1110101010110001),
    signed(1111010100110111),
    signed(1111100001000101),
    signed(1111011001010011),
    signed(0000010101100101),
    signed(1110110101010101),
    signed(1111001001011010),
    signed(1111011000011101),
    signed(1111010011100000),
    signed(1111101110100100),
    signed(1111010110011001),
    signed(0000100110110100),
    signed(0000011110011010),
    signed(0001100000011000),
    signed(0001001110101011),
    signed(0001010000011110),
    signed(0010100110000000),
    signed(0001101010010011),
    signed(0011101101001011),
    signed(0011010101110100),
    signed(0100100011011000),
    signed(0100111111101110),
    signed(0101010001001100),
    signed(0101101111010011),
    signed(0101101111111100),
    signed(0110110110101110),
    signed(0110101011011001),
    signed(0110001010100010),
    signed(0110010100000111),
    signed(0101111101110100),
    signed(0101110100111011),
    signed(0111101001111000),
    signed(0101011110001001),
    signed(0110101011001111),
    signed(0110001010111110),
    signed(0110101001001101),
    signed(0110000110011000),
    signed(0101100111111011),
    signed(0101010010111001),
    signed(0101100110000010),
    signed(0100101011101000),
    signed(0101100000010100),
    signed(0101001110010110),
    signed(0101010110110110),
    signed(0100110111011011),
    signed(0011101010111100),
    signed(0101000000110110),
    signed(0101001101110111),
    signed(0100001000010111),
    signed(0100101011000010),
    signed(0101100111100001),
    signed(0011101011111111),
    signed(0011010101100000),
    signed(0011110111010000),
    signed(0101001001100111),
    signed(0101010100101111),
    signed(0011101011111100),
    signed(0100000101101010),
    signed(0011110010010101),
    signed(0011110110100010),
    signed(0011011010100111),
    signed(0010110001011101),
    signed(0010111001101011),
    signed(0011000111100011),
    signed(0000101011111100),
    signed(0000110001110101),
    signed(0010011100100001),
    signed(1111101000110001),
    signed(1111110101101001),
    signed(1111011101001110),
    signed(1111000101110001),
    signed(1110100101101110),
    signed(1110000011010101),
    signed(1101101000111011),
    signed(1101111101110011),
    signed(1101010100010011),
    signed(1100111011110001),
    signed(1100101111011001),
    signed(1100110110000001),
    signed(1110000111111011),
    signed(1101010001010010),
    signed(1110010100001010),
    signed(1101100110100001),
    signed(1101101111011000),
    signed(1101101110011111),
    signed(1110010101000000),
    signed(1101111101111100),
    signed(1101110110111101),
    signed(1110001001101001),
    signed(1110101101000100),
    signed(1110011011100011),
    signed(1110111000111101),
    signed(1111010101000101),
    signed(0000000001101100),
    signed(1110010000100011),
    signed(1101100110111010),
    signed(1110010000100110),
    signed(1111000000101000),
    signed(1110000000001000),
    signed(1110011001101001),
    signed(1110000110010101),
    signed(1101100011011010),
    signed(1110010110100010),
    signed(1110011001110110),
    signed(1101111101001001),
    signed(1100111101011010),
    signed(1101100111000111),
    signed(1101000100010110),
    signed(1011111010001111),
    signed(1101011001111011),
    signed(1110011001001001),
    signed(1101001001110011),
    signed(1110100101111010),
    signed(1110111111111000),
    signed(1110000100101010),
    signed(1110010100001011),
    signed(1110011010110001),
    signed(1110110001011001),
    signed(1111001101001110),
    signed(1111011100101110),
    signed(1111000011100111),
    signed(1111101101111100),
    signed(0000010011011110),
    signed(0000111000111011),
    signed(0000000000110110),
    signed(1111001010110010),
    signed(1111011011001110),
    signed(1110101010001101),
    signed(1111100100000110),
    signed(1111111001001000),
    signed(1110100111001001),
    signed(1101100011011010),
    signed(1101010110000011),
    signed(1101110001100000),
    signed(1100101100110011),
    signed(1101010100101011),
    signed(1100100110001001),
    signed(1101011000110001),
    signed(1011110000101010),
    signed(1100000100100010),
    signed(1100110000010111),
    signed(1010101111101100),
    signed(1011010010011010),
    signed(1011000101010110),
    signed(1011100101000000),
    signed(1001101001111001),
    signed(1010000001101111),
    signed(1010010010101010),
    signed(1001101001101101),
    signed(1010100001011010),
    signed(1100000011100000),
    signed(1011010011001110),
    signed(1011100111000000),
    signed(1011000001100000),
    signed(1011111110110110),
    signed(1100110010010110),
    signed(1011101010000110),
    signed(1011101110111101),
    signed(1100111001000111),
    signed(1011010101011110),
    signed(1100110000111001),
    signed(1100000001101111),
    signed(1011111110001111),
    signed(1011101011110010),
    signed(1100001101100101),
    signed(1011111001101111),
    signed(1010101100010000),
    signed(1100110011010001),
    signed(1100001100011101),
    signed(1011000011111000),
    signed(1010101011010110),
    signed(1101001011011000),
    signed(1100010011111011),
    signed(1011010001110110),
    signed(1100010001001111),
    signed(1100011000011100),
    signed(1100010000011001),
    signed(1100110111011001),
    signed(1101101010100101),
    signed(1100110101100110),
    signed(1110101101011001),
    signed(1110100010011001),
    signed(1110111010111010),
    signed(1110111001001101),
);

begin
    
    data_out <= signal_array(to_integer(addr));

end Behaviroal;