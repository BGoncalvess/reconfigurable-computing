library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity filter_rom is
    Port ( 
        addr : in unsigned(5 downto 0);
        data_out : out signed(15 downto 0)
    );
end filter_rom;

architecture Behavioral of filter_rom is 

    type coeff_array is array (0 to 50) of signed(15 downto 0);

    constant coeffs : coeff_array := (
        "1111111110101011",
        "1111111110110001",
        "1111111110110011",
        "1111111110110101",
        "1111111110111001",
        "1111111111000100",
        "1111111111011000",
        "1111111111111010",
        "0000000000101011",
        "0000000001101111",
        "0000000011000110",
        "0000000100110000",
        "0000000110101101",
        "0000001000111011",
        "0000001011011000",
        "0000001101111111",
        "0000010000101101",
        "0000010011011101",
        "0000010110001010",
        "0000011000101101",
        "0000011011000010",
        "0000011101000100",
        "0000011110101110",
        "0000011111111100",
        "0000100000101100",
        "0000100000111101",
        "0000100000101100",
        "0000011111111100",
        "0000011110101110",
        "0000011101000100",
        "0000011011000010",
        "0000011000101101",
        "0000010110001010",
        "0000010011011101",
        "0000010000101101",
        "0000001101111111",
        "0000001011011000",
        "0000001000111011",
        "0000000110101101",
        "0000000100110000",
        "0000000011000110",
        "0000000001101111",
        "0000000000101011",
        "1111111111111010",
        "1111111111011000",
        "1111111111000100",
        "1111111110111001",
        "1111111110110101",
        "1111111110110011",
        "1111111110110001",
        "1111111110101011"
    );

begin
    data_out <= coeffs(to_integer(addr));
end Behavioral;
